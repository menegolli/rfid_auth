library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sine_mem is
	port (
		enable_mem		: std_logic;
		addr					: in std_logic_vector(7 downto 0);
		sine_mem_out 	: out std_logic_vector(7 downto 0)
	);
end entity sine_mem;

architecture sine_mem_arch of sine_mem is
	type mem is array ( 0 to 255 ) of std_logic_vector(7 downto 0);

	constant sine_samples : mem := (
		0    => "10000000",
		1    => "10000011",
		2    => "10000110",
		3    => "10001001",
		4    => "10001100",
		5    => "10001111",
		6    => "10010010",
		7    => "10010101",
		8    => "10011000",
		9    => "10011011",
		10   => "10011110",
		11   => "10100010",
		12   => "10100101",
		13   => "10100111",
		14   => "10101010",
		15   => "10101101",
		16   => "10110000",
		17   => "10110011",
		18   => "10110110",
		19   => "10111001",
		20   => "10111100",
		21   => "10111110",
		22   => "11000001",
		23   => "11000100",
		24   => "11000110",
		25   => "11001001",
		26   => "11001011",
		27   => "11001110",
		28   => "11010000",
		29   => "11010011",
		30   => "11010101",
		31   => "11010111",
		32   => "11011010",
		33   => "11011100",
		34   => "11011110",
		35   => "11100000",
		36   => "11100010",
		37   => "11100100",
		38   => "11100110",
		39   => "11101000",
		40   => "11101010",
		41   => "11101011",
		42   => "11101101",
		43   => "11101110",
		44   => "11110000",
		45   => "11110001",
		46   => "11110011",
		47   => "11110100",
		48   => "11110101",
		49   => "11110110",
		50   => "11111000",
		51   => "11111001",
		52   => "11111010",
		53   => "11111010",
		54   => "11111011",
		55   => "11111100",
		56   => "11111101",
		57   => "11111101",
		58   => "11111110",
		59   => "11111110",
		60   => "11111110",
		61   => "11111111",
		62   => "11111111",
		63   => "11111111",
		64   => "11111111",
		65   => "11111111",
		66   => "11111111",
		67   => "11111111",
		68   => "11111110",
		69   => "11111110",
		70   => "11111110",
		71   => "11111101",
		72   => "11111101",
		73   => "11111100",
		74   => "11111011",
		75   => "11111010",
		76   => "11111010",
		77   => "11111001",
		78   => "11111000",
		79   => "11110110",
		80   => "11110101",
		81   => "11110100",
		82   => "11110011",
		83   => "11110001",
		84   => "11110000",
		85   => "11101110",
		86   => "11101101",
		87   => "11101011",
		88   => "11101010",
		89   => "11101000",
		90   => "11100110",
		91   => "11100100",
		92   => "11100010",
		93   => "11100000",
		94   => "11011110",
		95   => "11011100",
		96   => "11011010",
		97   => "11010111",
		98   => "11010101",
		99   => "11010011",
		100  => "11010000",
		101  => "11001110",
		102  => "11001011",
		103  => "11001001",
		104  => "11000110",
		105  => "11000100",
		106  => "11000001",
		107  => "10111110",
		108  => "10111100",
		109  => "10111001",
		110  => "10110110",
		111  => "10110011",
		112  => "10110000",
		113  => "10101101",
		114  => "10101010",
		115  => "10100111",
		116  => "10100101",
		117  => "10100010",
		118  => "10011110",
		119  => "10011011",
		120  => "10011000",
		121  => "10010101",
		122  => "10010010",
		123  => "10001111",
		124  => "10001100",
		125  => "10001001",
		126  => "10000110",
		127  => "10000011",
		128  => "10000000",
		129  => "01111100",
		130  => "01111001",
		131  => "01110110",
		132  => "01110011",
		133  => "01110000",
		134  => "01101101",
		135  => "01101010",
		136  => "01100111",
		137  => "01100100",
		138  => "01100001",
		139  => "01011101",
		140  => "01011010",
		141  => "01011000",
		142  => "01010101",
		143  => "01010010",
		144  => "01001111",
		145  => "01001100",
		146  => "01001001",
		147  => "01000110",
		148  => "01000011",
		149  => "01000001",
		150  => "00111110",
		151  => "00111011",
		152  => "00111001",
		153  => "00110110",
		154  => "00110100",
		155  => "00110001",
		156  => "00101111",
		157  => "00101100",
		158  => "00101010",
		159  => "00101000",
		160  => "00100101",
		161  => "00100011",
		162  => "00100001",
		163  => "00011111",
		164  => "00011101",
		165  => "00011011",
		166  => "00011001",
		167  => "00010111",
		168  => "00010101",
		169  => "00010100",
		170  => "00010010",
		171  => "00010001",
		172  => "00001111",
		173  => "00001110",
		174  => "00001100",
		175  => "00001011",
		176  => "00001010",
		177  => "00001001",
		178  => "00000111",
		179  => "00000110",
		180  => "00000101",
		181  => "00000101",
		182  => "00000100",
		183  => "00000011",
		184  => "00000010",
		185  => "00000010",
		186  => "00000001",
		187  => "00000001",
		188  => "00000001",
		189  => "00000000",
		190  => "00000000",
		191  => "00000000",
		192  => "00000000",
		193  => "00000000",
		194  => "00000000",
		195  => "00000000",
		196  => "00000001",
		197  => "00000001",
		198  => "00000001",
		199  => "00000010",
		200  => "00000010",
		201  => "00000011",
		202  => "00000100",
		203  => "00000101",
		204  => "00000101",
		205  => "00000110",
		206  => "00000111",
		207  => "00001001",
		208  => "00001010",
		209  => "00001011",
		210  => "00001100",
		211  => "00001110",
		212  => "00001111",
		213  => "00010001",
		214  => "00010010",
		215  => "00010100",
		216  => "00010101",
		217  => "00010111",
		218  => "00011001",
		219  => "00011011",
		220  => "00011101",
		221  => "00011111",
		222  => "00100001",
		223  => "00100011",
		224  => "00100101",
		225  => "00101000",
		226  => "00101010",
		227  => "00101100",
		228  => "00101111",
		229  => "00110001",
		230  => "00110100",
		231  => "00110110",
		232  => "00111001",
		233  => "00111011",
		234  => "00111110",
		235  => "01000001",
		236  => "01000011",
		237  => "01000110",
		238  => "01001001",
		239  => "01001100",
		240  => "01001111",
		241  => "01010010",
		242  => "01010101",
		243  => "01011000",
		244  => "01011010",
		245  => "01011101",
		246  => "01100001",
		247  => "01100100",
		248  => "01100111",
		249  => "01101010",
		250  => "01101101",
		251  => "01110000",
		252  => "01110011",
		253  => "01110110",
		254  => "01111001",
		255  => "01111100"
	);

begin
	mem_out : process(enable_mem, addr)
	begin
		if enable_mem = '1' then
			sine_mem_out <= sine_samples(to_integer(unsigned(addr)));
		else
			sine_mem_out <= (others => '0');
		end if;
	end process;
end architecture sine_mem_arch;
